package mypkg;
	 import   uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "my_config.svh"
	`include "my_transaction.svh"
	`include "my_driver.svh"
	`include "my_sequencer.svh"
	`include "my_agent.svh"
	//`include "my_env.svh"
	//`include "my_test.svh"
endpackage